
package env_defines;
typedef enum {ADDR_7_BIT,ADDR_10_BIT} slave_addr_mode;
typedef enum {FREE,BUSY} bfm_stat;
endpackage

